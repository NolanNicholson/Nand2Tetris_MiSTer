// gate names are reserved identifiers in Verilog; hence the "_n2t" suffix
module not_n2t
(
    input in,
    output out
);

// TODO

endmodule
