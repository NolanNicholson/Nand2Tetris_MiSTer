module Add16
(
    input [15:0] a,
    input [15:0] b,

    output [15:0] out
);

// TODO

endmodule
