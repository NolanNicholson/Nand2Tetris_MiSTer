// DESCRIPTION: Verilator: Verilog example module
//
// This file ONLY is placed under the Creative Commons Public Domain, for
// any use, without warranty, 2017 by Wilson Snyder.
// SPDX-License-Identifier: CC0-1.0

// See also https://verilator.org/guide/latest/examples.html"

module top
(
    input in_a,
    input in_b,
    output out_nand
);

nand_n2t nand01
(
    .a(in_a),
    .b(in_b),
    .out(out_nand)
);

endmodule
