module HackALU
(
    input [15:0] x,
    input [15:0] y,

    output [15:0] out,

    input zx,
    input nx,
    input zy,
    input ny,
    input f,
    input no,

    output zr,
    output ng
);

// TODO

endmodule
