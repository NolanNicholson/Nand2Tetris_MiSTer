module dmux4way
(
    input in,
    input [1:0] sel,
    output a,
    output b,
    output c,
    output d
);

// TODO

endmodule
