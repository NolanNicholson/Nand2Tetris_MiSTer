// gate names are reserved identifiers in Verilog; hence the "_n2t" suffix
module xor_n2t
(
    input a,
    input b,
    output out
);

// TODO

endmodule
