module and16
(
    input [15:0] a,
    input [15:0] b,
    output [15:0] out
);


and_n2t and0
(
    .a(a[0]),
    .b(b[0]),
    .out(out[0])
);

and_n2t and1
(
    .a(a[1]),
    .b(b[1]),
    .out(out[1])
);

and_n2t and2
(
    .a(a[2]),
    .b(b[2]),
    .out(out[2])
);

and_n2t and3
(
    .a(a[3]),
    .b(b[3]),
    .out(out[3])
);

and_n2t and4
(
    .a(a[4]),
    .b(b[4]),
    .out(out[4])
);

and_n2t and5
(
    .a(a[5]),
    .b(b[5]),
    .out(out[5])
);

and_n2t and6
(
    .a(a[6]),
    .b(b[6]),
    .out(out[6])
);

and_n2t and7
(
    .a(a[7]),
    .b(b[7]),
    .out(out[7])
);

and_n2t and8
(
    .a(a[8]),
    .b(b[8]),
    .out(out[8])
);

and_n2t and9
(
    .a(a[9]),
    .b(b[9]),
    .out(out[9])
);

and_n2t and10
(
    .a(a[10]),
    .b(b[10]),
    .out(out[10])
);

and_n2t and11
(
    .a(a[11]),
    .b(b[11]),
    .out(out[11])
);

and_n2t and12
(
    .a(a[12]),
    .b(b[12]),
    .out(out[12])
);

and_n2t and13
(
    .a(a[13]),
    .b(b[13]),
    .out(out[13])
);

and_n2t and14
(
    .a(a[14]),
    .b(b[14]),
    .out(out[14])
);

and_n2t and15
(
    .a(a[15]),
    .b(b[15]),
    .out(out[15])
);


endmodule
