module dmux
(
    input in,
    input sel,
    output a,
    output b
);

// TODO

endmodule
