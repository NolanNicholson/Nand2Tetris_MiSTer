module FullAdder
(
    input a,
    input b,
    input c,
    output sum,
    output carry
);

// TODO

endmodule
