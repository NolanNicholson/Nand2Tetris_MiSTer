module mux
(
    input a,
    input b,
    input sel,
    output out
);

// TODO

endmodule
