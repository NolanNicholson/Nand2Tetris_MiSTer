module or8way
(
    input [7:0] in,
    output out
);

// TODO

endmodule
