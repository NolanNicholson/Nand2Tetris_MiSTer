module Inc16
(
    input [15:0] in,
    output [15:0] out
);

// TODO

endmodule
